library ieee;
use ieee.std_logic_1164.all;

entity map4 is
	port
	(
		F0, F1, F2, F3, F4, F5, F6, F7, F8, F9, F10, F11, F12, F13, F14, F15: out std_logic_vector(31 downto 0)
	);
end map4;	
	
architecture map4_struct of map4 is
begin
	F0 <=  "11111111111111111111111111111111";
	F1 <=  "00110000000001111110000000001110";
	F2 <=  "00000000000000000001110000000000";
	F3 <=  "00000000111110000000000000000000";
	F4 <=  "00000000000000001110000000111000";
	F5 <=  "01100000000000000000000000001111";
	F6 <=  "00000000011111100000001110000000";
	F7 <=  "00000000000000000111000000000000";
	F8 <=  "00111000000000111111111111111111";
	F9 <=  "01110000000000111111111100100010";
	F10<=  "00000001111111111111000000001010";
	F11<=  "00000000001000000000000100000000";
	F12<=  "00011111000011000001000001000010";
	F13<=  "00111110011000001100001000000000";
	F14<=  "01111100000001111100000000010000";
	F15<=  "11111111111111111111111111111111";
end map4_struct;