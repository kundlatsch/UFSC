library ieee;
use ieee.std_logic_1164.all;

entity map3 is
	port
	(
		F0, F1, F2, F3, F4, F5, F6, F7, F8, F9, F10, F11, F12, F13, F14, F15: out std_logic_vector(31 downto 0)
	);
end map3;	
	
architecture map3_struct of map3 is
begin
	F0 <=  "00000000011111111111000000000000";
	F1 <=  "00000000000000011111111111110000";
	F2 <=  "00000011111100000000000000000000";
	F3 <=  "00000111111111111000000100010000";
	F4 <=  "00010000011000000000000000000000";
	F5 <=  "00000000001100110110011000000111";
	F6 <=  "00000000001110000000000000000000";
	F7 <=  "00000000011111111110000000000000";
	F8 <=  "00000000000000000000000000000000";
	F9 <=  "00000000001000000111100000100000";
	F10<=  "00010000010000011100000000000000";
	F11<=  "00000000000010010000000000001000";
	F12<=  "00000000000011110000000000100000";
	F13<=  "00100001111110000000011110000000";
	F14<=  "00000000000000001110000000000000";
	F15<=  "00010000011111111111110000000100";
end map3_struct;